<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-4.83236,-3.87211,104.09,-57.7106</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>34.5,-8</position>
<gparam>LABEL_TEXT Design 4X16 decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>BI_DECODER_4x16</type>
<position>29,-24.5</position>
<input>
<ID>ENABLE</ID>5 </input>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_10</ID>15 </output>
<output>
<ID>OUT_11</ID>14 </output>
<output>
<ID>OUT_12</ID>12 </output>
<output>
<ID>OUT_13</ID>10 </output>
<output>
<ID>OUT_14</ID>3 </output>
<output>
<ID>OUT_15</ID>2 </output>
<output>
<ID>OUT_2</ID>23 </output>
<output>
<ID>OUT_3</ID>22 </output>
<output>
<ID>OUT_4</ID>21 </output>
<output>
<ID>OUT_5</ID>20 </output>
<output>
<ID>OUT_6</ID>19 </output>
<output>
<ID>OUT_7</ID>18 </output>
<output>
<ID>OUT_8</ID>17 </output>
<output>
<ID>OUT_9</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>36.5,-11</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>36.5,-13.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>36.5,-16</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>36.5,-18.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>36.5,-36</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>36.5,-21</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>36.5,-23.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>36.5,-31</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>36.5,-26</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>36.5,-38.5</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>36.5,-33.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>36.5,-28.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>36.5,-41</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>36.5,-43.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>36.5,-48.5</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>36.5,-46</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>22.5,-15</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>21,-25</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>21,-27.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>21,-30</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>21,-32.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>61,-24</position>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-17,33.5,-11</points>
<intersection>-17 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-11,35.5,-11</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-17,33.5,-17</points>
<connection>
<GID>4</GID>
<name>OUT_15</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-13.5,35.5,-13.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>34 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>34,-18,34,-13.5</points>
<intersection>-18 5</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>32,-18,34,-18</points>
<connection>
<GID>4</GID>
<name>OUT_14</name></connection>
<intersection>34 4</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-17,25.5,-15</points>
<intersection>-17 3</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-15,25.5,-15</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-17,26,-17</points>
<connection>
<GID>4</GID>
<name>ENABLE</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-29,25,-25</points>
<intersection>-29 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-29,26,-29</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-25,25,-25</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-30,25,-27.5</points>
<intersection>-30 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-30,26,-30</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-27.5,25,-27.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-31,24.5,-30</points>
<intersection>-31 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-31,26,-31</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-30,24.5,-30</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-32.5,24.5,-32</points>
<intersection>-32.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-32,26,-32</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-32.5,24.5,-32.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-19,33.5,-16</points>
<intersection>-19 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-16,35.5,-16</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-19,33.5,-19</points>
<connection>
<GID>4</GID>
<name>OUT_13</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-20,35.5,-20</points>
<connection>
<GID>4</GID>
<name>OUT_12</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-20,35.5,-18.5</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-21,35.5,-21</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-22,35.5,-22</points>
<connection>
<GID>4</GID>
<name>OUT_10</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-23.5,35.5,-22</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-26,34,-23</points>
<intersection>-26 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-26,35.5,-26</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-23,34,-23</points>
<connection>
<GID>4</GID>
<name>OUT_9</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-28.5,34,-24</points>
<intersection>-28.5 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-28.5,35.5,-28.5</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-24,34,-24</points>
<connection>
<GID>4</GID>
<name>OUT_8</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-31,34,-25</points>
<intersection>-31 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-31,35.5,-31</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-25,34,-25</points>
<connection>
<GID>4</GID>
<name>OUT_7</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-33.5,34,-26</points>
<intersection>-33.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-33.5,35.5,-33.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-26,34,-26</points>
<connection>
<GID>4</GID>
<name>OUT_6</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-36,34,-27</points>
<intersection>-36 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-36,35.5,-36</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-27,34,-27</points>
<connection>
<GID>4</GID>
<name>OUT_5</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-38.5,34,-28</points>
<intersection>-38.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-38.5,35.5,-38.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-28,34,-28</points>
<connection>
<GID>4</GID>
<name>OUT_4</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-41,34,-29</points>
<intersection>-41 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-41,35.5,-41</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-29,34,-29</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-43.5,34,-30</points>
<intersection>-43.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-43.5,35.5,-43.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-30,34,-30</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-46,33.5,-31</points>
<intersection>-46 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-46,35.5,-46</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-31,33.5,-31</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-48.5,33.5,-32</points>
<intersection>-48.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-48.5,35.5,-48.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-32,33.5,-32</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-14.9208,13.3065,199.75,-92.8014</PageViewport>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>37,-4.5</position>
<gparam>LABEL_TEXT 4X16 using 3X8 Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>BE_DECODER_3x8</type>
<position>26,-18.5</position>
<input>
<ID>ENABLE</ID>29 </input>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT_0</ID>38 </output>
<output>
<ID>OUT_1</ID>37 </output>
<output>
<ID>OUT_2</ID>36 </output>
<output>
<ID>OUT_3</ID>35 </output>
<output>
<ID>OUT_4</ID>34 </output>
<output>
<ID>OUT_5</ID>33 </output>
<output>
<ID>OUT_6</ID>32 </output>
<output>
<ID>OUT_7</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>60</ID>
<type>BE_DECODER_3x8</type>
<position>25.5,-42</position>
<input>
<ID>ENABLE</ID>30 </input>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT_0</ID>48 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_2</ID>46 </output>
<output>
<ID>OUT_3</ID>45 </output>
<output>
<ID>OUT_4</ID>44 </output>
<output>
<ID>OUT_5</ID>42 </output>
<output>
<ID>OUT_6</ID>41 </output>
<output>
<ID>OUT_7</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>3,-18.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>4,-22</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>3,-15.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>5.5,-10</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_INVERTER</type>
<position>14.5,-8.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>31.5,-11.5</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>31.5,-14</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>31.5,-16.5</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>31.5,-19</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>31.5,-21.5</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>31.5,-24</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>31.5,-9</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>31.5,-26.5</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>31.5,-36.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>31.5,-39</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>31.5,-41.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>31.5,-44</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>GA_LED</type>
<position>31.5,-46.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>31.5,-49</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>31.5,-34</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>31.5,-51.5</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-20,11,-15.5</points>
<intersection>-20 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-20,23,-20</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>11 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-15.5,11,-15.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-43.5,15.5,-20</points>
<intersection>-43.5 4</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-43.5,22.5,-43.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-21,11,-18.5</points>
<intersection>-21 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-21,23,-21</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection>
<intersection>14.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-18.5,11,-18.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-44.5,14.5,-21</points>
<intersection>-44.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-44.5,22.5,-44.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-22,23,-22</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>16.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-45.5,16.5,-22</points>
<intersection>-45.5 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16.5,-45.5,22.5,-45.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>16.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-15,10.5,-8.5</points>
<intersection>-15 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-15,23,-15</points>
<connection>
<GID>58</GID>
<name>ENABLE</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-8.5,11.5,-8.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>7.5 4</intersection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>7.5,-10,7.5,-8.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-38.5,20,-8.5</points>
<intersection>-38.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-38.5,22.5,-38.5</points>
<connection>
<GID>60</GID>
<name>ENABLE</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-8.5,20,-8.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-15,29.5,-9</points>
<intersection>-15 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-9,30.5,-9</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-15,29.5,-15</points>
<connection>
<GID>58</GID>
<name>OUT_7</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-16,29.5,-11.5</points>
<intersection>-16 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-11.5,30.5,-11.5</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-16,29.5,-16</points>
<connection>
<GID>58</GID>
<name>OUT_6</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-17,29.5,-14</points>
<intersection>-17 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-14,30.5,-14</points>
<connection>
<GID>74</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-17,29.5,-17</points>
<connection>
<GID>58</GID>
<name>OUT_5</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-18,29.5,-16.5</points>
<intersection>-18 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-16.5,30.5,-16.5</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-18,29.5,-18</points>
<connection>
<GID>58</GID>
<name>OUT_4</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-19,30.5,-19</points>
<connection>
<GID>78</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-21.5,29.5,-20</points>
<intersection>-21.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-21.5,30.5,-21.5</points>
<connection>
<GID>80</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-20,29.5,-20</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-24,29.5,-21</points>
<intersection>-24 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-24,30.5,-24</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-21,29.5,-21</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-26.5,29.5,-22</points>
<intersection>-26.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-26.5,30.5,-26.5</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-22,29.5,-22</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-38.5,29,-34</points>
<intersection>-38.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-34,30.5,-34</points>
<connection>
<GID>93</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-38.5,29,-38.5</points>
<connection>
<GID>60</GID>
<name>OUT_7</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-39.5,29,-36.5</points>
<intersection>-39.5 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-36.5,30.5,-36.5</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-39.5,29,-39.5</points>
<connection>
<GID>60</GID>
<name>OUT_6</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-40.5,29,-39</points>
<intersection>-40.5 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-39,30.5,-39</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-40.5,29,-40.5</points>
<connection>
<GID>60</GID>
<name>OUT_5</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-41.5,30.5,-41.5</points>
<connection>
<GID>60</GID>
<name>OUT_4</name></connection>
<connection>
<GID>89</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-44,29,-42.5</points>
<intersection>-44 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-44,30.5,-44</points>
<connection>
<GID>90</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-42.5,29,-42.5</points>
<connection>
<GID>60</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-46.5,29,-43.5</points>
<intersection>-46.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-46.5,30.5,-46.5</points>
<connection>
<GID>91</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-43.5,29,-43.5</points>
<connection>
<GID>60</GID>
<name>OUT_2</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-49,29,-44.5</points>
<intersection>-49 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-49,30.5,-49</points>
<connection>
<GID>92</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-44.5,29,-44.5</points>
<connection>
<GID>60</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-51.5,29,-45.5</points>
<intersection>-51.5 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-51.5,30.5,-51.5</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-45.5,29,-45.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-47.5076,2.09721,74.8924,-58.4028</PageViewport>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>20.5,-8</position>
<gparam>LABEL_TEXT 4X16 using 2X4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>BA_DECODER_2x4</type>
<position>22.5,-19.5</position>
<input>
<ID>ENABLE</ID>49 </input>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT_0</ID>65 </output>
<output>
<ID>OUT_1</ID>62 </output>
<output>
<ID>OUT_2</ID>63 </output>
<output>
<ID>OUT_3</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>BA_DECODER_2x4</type>
<position>23,-28.5</position>
<input>
<ID>ENABLE</ID>50 </input>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT_0</ID>69 </output>
<output>
<ID>OUT_1</ID>68 </output>
<output>
<ID>OUT_2</ID>67 </output>
<output>
<ID>OUT_3</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>BA_DECODER_2x4</type>
<position>23,-37</position>
<input>
<ID>ENABLE</ID>55 </input>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT_0</ID>73 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>71 </output>
<output>
<ID>OUT_3</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_DECODER_2x4</type>
<position>23.5,-46.5</position>
<input>
<ID>ENABLE</ID>52 </input>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT_0</ID>77 </output>
<output>
<ID>OUT_1</ID>76 </output>
<output>
<ID>OUT_2</ID>75 </output>
<output>
<ID>OUT_3</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>BA_DECODER_2x4</type>
<position>-5,-30.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT_0</ID>52 </output>
<output>
<ID>OUT_1</ID>55 </output>
<output>
<ID>OUT_2</ID>50 </output>
<output>
<ID>OUT_3</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>-12,-31</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>-12,-35</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-15.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-18.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>33.5,-11.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>33.5,-14</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>33.5,-16.5</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>33.5,-19</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>GA_LED</type>
<position>33.5,-22.5</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>33.5,-25</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>33.5,-27.5</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>GA_LED</type>
<position>33.5,-30</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>33.5,-33</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>GA_LED</type>
<position>33.5,-35.5</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>GA_LED</type>
<position>33.5,-38</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>33.5,-40.5</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>GA_LED</type>
<position>33.5,-44</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>33.5,-46.5</position>
<input>
<ID>N_in0</ID>75 </input>
<input>
<ID>N_in1</ID>78 </input>
<input>
<ID>N_in3</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>33.5,-49</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>33.5,-51.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-29,6,-18</points>
<intersection>-29 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-18,19.5,-18</points>
<connection>
<GID>100</GID>
<name>ENABLE</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-29,6,-29</points>
<connection>
<GID>108</GID>
<name>OUT_3</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-30,6,-29</points>
<intersection>-30 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-29,20,-29</points>
<intersection>6 0</intersection>
<intersection>20 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-30,6,-30</points>
<connection>
<GID>108</GID>
<name>OUT_2</name></connection>
<intersection>6 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-29,20,-27</points>
<connection>
<GID>102</GID>
<name>ENABLE</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-45,5,-32</points>
<intersection>-45 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-45,20.5,-45</points>
<connection>
<GID>106</GID>
<name>ENABLE</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-32,5,-32</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-35,-8.5,-32</points>
<intersection>-35 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-32,-8,-32</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-35,-8.5,-35</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-31,-8,-31</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-35.5,6,-31</points>
<intersection>-35.5 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-35.5,20,-35.5</points>
<connection>
<GID>104</GID>
<name>ENABLE</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-31,6,-31</points>
<connection>
<GID>108</GID>
<name>OUT_1</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-21,0.5,-18.5</points>
<intersection>-21 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-21,19.5,-21</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-18.5,0.5,-18.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-48,15.5,-21</points>
<intersection>-48 8</intersection>
<intersection>-38.5 7</intersection>
<intersection>-30 6</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>15.5,-30,20,-30</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>15.5,-38.5,20,-38.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>15.5,-48,20.5,-48</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-15.5,19.5,-15.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>14 3</intersection>
<intersection>19.5 14</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-47,14,-15.5</points>
<intersection>-47 12</intersection>
<intersection>-37.5 10</intersection>
<intersection>-29 9</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>14,-29,20,-29</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>14 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14,-37.5,20,-37.5</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>14 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>14,-47,20.5,-47</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>14 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>19.5,-20,19.5,-15.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-20,26,-16.5</points>
<intersection>-20 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-16.5,32.5,-16.5</points>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-20,26,-20</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-19,26,-14</points>
<intersection>-19 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-14,32.5,-14</points>
<connection>
<GID>122</GID>
<name>N_in0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-19,26,-19</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-18,26,-11.5</points>
<intersection>-18 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-11.5,32.5,-11.5</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-18,26,-18</points>
<connection>
<GID>100</GID>
<name>OUT_3</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-21,26,-19</points>
<intersection>-21 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-19,32.5,-19</points>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-21,26,-21</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-27,29,-22.5</points>
<intersection>-27 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-22.5,32.5,-22.5</points>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-27,29,-27</points>
<connection>
<GID>102</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-28,29,-25</points>
<intersection>-28 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-25,32.5,-25</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-28,29,-28</points>
<connection>
<GID>102</GID>
<name>OUT_2</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-29,29,-27.5</points>
<intersection>-29 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-27.5,32.5,-27.5</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-29,29,-29</points>
<connection>
<GID>102</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-30,32.5,-30</points>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-35.5,29,-33</points>
<intersection>-35.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-33,32.5,-33</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-35.5,29,-35.5</points>
<connection>
<GID>104</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-36.5,29,-35.5</points>
<intersection>-36.5 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-35.5,32.5,-35.5</points>
<connection>
<GID>132</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-36.5,29,-36.5</points>
<connection>
<GID>104</GID>
<name>OUT_2</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-38,29,-37.5</points>
<intersection>-38 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-38,32.5,-38</points>
<connection>
<GID>133</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-37.5,29,-37.5</points>
<connection>
<GID>104</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-40.5,29,-38.5</points>
<intersection>-40.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-40.5,32.5,-40.5</points>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-38.5,29,-38.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-45,29.5,-44</points>
<intersection>-45 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-44,32.5,-44</points>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-45,29.5,-45</points>
<connection>
<GID>106</GID>
<name>OUT_3</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-46.5,29.5,-46</points>
<intersection>-46.5 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-46.5,32.5,-46.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-46,29.5,-46</points>
<connection>
<GID>106</GID>
<name>OUT_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-49,33.5,-48</points>
<connection>
<GID>137</GID>
<name>N_in3</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-49,33.5,-49</points>
<intersection>30 2</intersection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>30,-49,30,-47</points>
<intersection>-49 1</intersection>
<intersection>-47 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-47,30,-47</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<intersection>30 2</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-51.5,29.5,-48</points>
<intersection>-51.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-51.5,32.5,-51.5</points>
<connection>
<GID>138</GID>
<name>N_in0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-48,29.5,-48</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-46,33.5,-45.5</points>
<connection>
<GID>136</GID>
<name>N_in3</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-46,34.5,-46</points>
<intersection>33.5 0</intersection>
<intersection>34.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>34.5,-46.5,34.5,-46</points>
<connection>
<GID>136</GID>
<name>N_in1</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-0.594141,-8.74766,57.498,-37.4615</PageViewport>
<gate>
<ID>144</ID>
<type>AE_DFF_LOW</type>
<position>41,-16</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUTINV_0</ID>90 </output>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>148</ID>
<type>BB_CLOCK</type>
<position>12,-19.5</position>
<output>
<ID>CLK</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>21.5,-21.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>152</ID>
<type>DA_FROM</type>
<position>30.5,-17</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>30,-14</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>156</ID>
<type>DE_TO</type>
<position>26,-12</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_TOGGLE</type>
<position>20.5,-12</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>3.5,-16</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>47.5,-14</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q</lparam></gate>
<gate>
<ID>164</ID>
<type>GA_LED</type>
<position>8,-16</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>3.5,-20</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q'</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>46.5,-17</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q'</lparam></gate>
<gate>
<ID>170</ID>
<type>GA_LED</type>
<position>6.5,-20</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-21.5,17.5,-19.5</points>
<intersection>-21.5 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-21.5,19.5,-21.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-19.5,17.5,-19.5</points>
<connection>
<GID>148</GID>
<name>CLK</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-17,38,-17</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-12,24,-12</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>22.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22.5,-12,22.5,-12</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-14,38,-14</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-14,45.5,-14</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-14,44,-14</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-16,7,-16</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>7 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7,-16,7,-16</points>
<connection>
<GID>164</GID>
<name>N_in0</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-17,44.5,-17</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>44 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>44,-17,44,-17</points>
<connection>
<GID>144</GID>
<name>OUTINV_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-20,5.5,-20</points>
<connection>
<GID>170</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>