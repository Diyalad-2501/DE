<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>16.844,-10.4328,162.644,-84.1328</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>31.5,-19.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>23.5,-18</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>24,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>37.5,-19.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>31,-13</position>
<gparam>LABEL_TEXT AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR2</type>
<position>65,-20</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>58.5,-18</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>58.5,-22</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>69,-20</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>64.5,-13</position>
<gparam>LABEL_TEXT OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>BA_NAND2</type>
<position>31.5,-36</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>25.5,-34</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>25,-37.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AI_XOR2</type>
<position>63,-35</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>56.5,-33</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>56.5,-37</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>67,-35</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>63,-28</position>
<gparam>LABEL_TEXT XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>30.5,-29.5</position>
<gparam>LABEL_TEXT NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>40,-36</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-18.5,28.5,-18.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-18.5,26,-18</points>
<intersection>-18.5 1</intersection>
<intersection>-18 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-18,26,-18</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>26 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-21.5,27,-20.5</points>
<intersection>-21.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-21.5,27,-21.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-20.5,28.5,-20.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>34.5,-19.5,36.5,-19.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-19,62,-18</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-18,62,-18</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-22,62,-21</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-22,62,-22</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-20,68,-20</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-34,28.5,-34</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-35,28.5,-34</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-34,60,-33</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-33,60,-33</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-35,66,-35</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-37,60,-36</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-37,60,-37</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-36,39,-36</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-37.5,28,-37</points>
<intersection>-37.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-37,28.5,-37</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-37.5,28,-37.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-8.56149,7.24699,137.239,-66.453</PageViewport>
<gate>
<ID>42</ID>
<type>BA_NAND2</type>
<position>13,-15</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>3.5,-14</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>22.5,-15</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>16,-9.5</position>
<gparam>LABEL_TEXT NOT using NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>60.5,-1.5</position>
<gparam>LABEL_TEXT NAND as Universal Gate</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>14,-27.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>8,-25.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>8,-30</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>-62,-12.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>23,-27.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>29,-27.5</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>BA_NAND2</type>
<position>58,-27</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_NAND2</type>
<position>58,-32.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>51,-25.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>51.5,-34</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>BA_NAND2</type>
<position>67.5,-29</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>74.5,-29</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>16,-22</position>
<gparam>LABEL_TEXT AND using NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>64.5,-21.5</position>
<gparam>LABEL_TEXT OR using NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-16,7,-14</points>
<intersection>-16 3</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-14,10,-14</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>7,-16,10,-16</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-15,21.5,-15</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-26.5,11,-25.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-25.5,11,-25.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-30,11,-28.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-30 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>10,-30,11,-30</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-27.5,28,-27.5</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-28.5,18.5,-26.5</points>
<intersection>-28.5 3</intersection>
<intersection>-27.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-26.5,20,-26.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-27.5,18.5,-27.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>18.5,-28.5,20,-28.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-28,55,-25.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-25.5,55,-25.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-34,55,-31.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-34,55,-34</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-28,62.5,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-28,64.5,-28</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-27,62.5,-27</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-32.5,62.5,-30</points>
<intersection>-32.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-30,64.5,-30</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-32.5,62.5,-32.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-29,73.5,-29</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<connection>
<GID>88</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>47.5,-3.5</position>
<gparam>LABEL_TEXT X-OR using NOR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>BE_NOR2</type>
<position>20,-18.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>BE_NOR2</type>
<position>21,-32</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>15,-17.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>14,-33</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>12.5,-17.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>12,-33</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>BE_NOR2</type>
<position>32,-21.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>BE_NOR2</type>
<position>33.5,-30</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>BE_NOR2</type>
<position>42,-25.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>BE_NOR2</type>
<position>52,-25</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>58,-25</position>
<input>
<ID>N_in2</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-25,17,-17.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-25,29.5,-25</points>
<intersection>17 0</intersection>
<intersection>29.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>29.5,-29,29.5,-25</points>
<intersection>-29 3</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-29,30.5,-29</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-33,18,-33</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>18 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>18,-33,18,-22.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>-33 1</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>18,-22.5,29,-22.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>18 4</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-20.5,26,-18.5</points>
<intersection>-20.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-20.5,29,-20.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-18.5,26,-18.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-32,26.5,-31</points>
<intersection>-32 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-31,30.5,-31</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-32,26.5,-32</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-24.5,37,-21.5</points>
<intersection>-24.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-24.5,39,-24.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-21.5,37,-21.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-30,37.5,-26.5</points>
<intersection>-30 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-26.5,39,-26.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-30,37.5,-30</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-25.5,47,-24</points>
<intersection>-25.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-24,49,-24</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection>
<intersection>49 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-25.5,47,-25.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-26,49,-24</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-26,58,-25</points>
<connection>
<GID>118</GID>
<name>N_in2</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-25,58,-25</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport>
<gate>
<ID>122</ID>
<type>AA_AND3</type>
<position>55.5,-26</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>32,-24</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>32,-30</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>32,-34.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_INVERTER</type>
<position>41,-29</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND2</type>
<position>55.5,-36.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_OR2</type>
<position>65,-31</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>72.5,-31</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>53.5,-4</position>
<gparam>LABEL_TEXT y=AB'C+B'C</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-35.5,47,-26</points>
<intersection>-35.5 9</intersection>
<intersection>-29 8</intersection>
<intersection>-26 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>44,-29,47,-29</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>47,-35.5,52.5,-35.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>47,-26,52.5,-26</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-29,38,-29</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>34 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>34,-30,34,-29</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-24,52.5,-24</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-37.5,45,-28</points>
<intersection>-37.5 3</intersection>
<intersection>-34.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-28,52.5,-28</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-34.5,45,-34.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45,-37.5,52.5,-37.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-30,59,-26</points>
<intersection>-30 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-30,62,-30</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-26,59,-26</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-36.5,59,-32</points>
<intersection>-36.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-32,62,-32</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-36.5,59,-36.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-31,71.5,-31</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<connection>
<GID>136</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-18,0,127.8,-73.7</PageViewport>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>63.5,-4.5</position>
<gparam>LABEL_TEXT Half Adder using NAND Gate</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>BA_NAND2</type>
<position>18.5,-17</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>BA_NAND2</type>
<position>18.5,-25</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>11,-15.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>11.5,-27</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>9,-15</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>9,-27</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BE_NOR2</type>
<position>-52,-29.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>BA_NAND2</type>
<position>29.5,-17</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>BA_NAND2</type>
<position>31,-26.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>BA_NAND2</type>
<position>41,-21</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>47.5,-21</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>BA_NAND2</type>
<position>27.5,-35</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>BA_NAND2</type>
<position>37,-35</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>GA_LED</type>
<position>43,-34.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-15.5,15.5,-15.5</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>15 5</intersection>
<intersection>15.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-18,15.5,-15.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>15,-34,15,-15.5</points>
<intersection>-34 6</intersection>
<intersection>-16 7</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>15,-34,24.5,-34</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>15 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>15,-16,26.5,-16</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>15 5</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-36,14.5,-27.5</points>
<intersection>-36 8</intersection>
<intersection>-29 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-29,28,-29</points>
<intersection>14.5 0</intersection>
<intersection>15.5 3</intersection>
<intersection>28 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-27.5,14.5,-27.5</points>
<intersection>14 4</intersection>
<intersection>14.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-29,15.5,-24</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>-29 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>14,-27.5,14,-27</points>
<intersection>-27.5 2</intersection>
<intersection>-27 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>13.5,-27,14,-27</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>14 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>28,-29,28,-27.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>14.5,-36,24.5,-36</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-25,24,-18</points>
<intersection>-25 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-18,26.5,-18</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-25,24,-25</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-25.5,24.5,-17</points>
<intersection>-25.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-25.5,28,-25.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-17,24.5,-17</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-20,35,-17</points>
<intersection>-20 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-20,38,-20</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-17,35,-17</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-26.5,36,-22</points>
<intersection>-26.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-22,38,-22</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-26.5,36,-26.5</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-35,34,-35</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-36,34,-34</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-35,41,-34.5</points>
<intersection>-35 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-34.5,42,-34.5</points>
<connection>
<GID>168</GID>
<name>N_in0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-35,41,-35</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-21,46.5,-21</points>
<connection>
<GID>162</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport>
<gate>
<ID>194</ID>
<type>AA_AND3</type>
<position>43.5,-18.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND3</type>
<position>43.5,-28</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>72 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND3</type>
<position>47,-38.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>72 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND3</type>
<position>44.5,-47</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_OR4</type>
<position>58,-27.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<input>
<ID>IN_2</ID>75 </input>
<input>
<ID>IN_3</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>204</ID>
<type>GA_LED</type>
<position>64.5,-27.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AE_OR3</type>
<position>59.5,-61.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<input>
<ID>IN_2</ID>80 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND2</type>
<position>47,-56</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>45,-63.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>45,-70.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>GA_LED</type>
<position>64.5,-62</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>52.5,-3.5</position>
<gparam>LABEL_TEXT Full Subtractor using AOI</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_INVERTER</type>
<position>24,-19</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_INVERTER</type>
<position>23.5,-25.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_TOGGLE</type>
<position>4.5,-21</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>4.5,-28</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>4.5,-35</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_INVERTER</type>
<position>26.5,-33</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-52.5,38.5,-52.5</points>
<intersection>15 14</intersection>
<intersection>21 15</intersection>
<intersection>38.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>38.5,-52.5,38.5,-36.5</points>
<intersection>-52.5 1</intersection>
<intersection>-45 9</intersection>
<intersection>-36.5 13</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>38.5,-45,41.5,-45</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>38.5 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>38.5,-36.5,44,-36.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>38.5 8</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>15,-52.5,15,-21</points>
<intersection>-52.5 1</intersection>
<intersection>-21 16</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>21,-52.5,21,-19</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>6.5,-21,15,-21</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>15 14</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-30,30.5,-30</points>
<intersection>16.5 5</intersection>
<intersection>21 6</intersection>
<intersection>24 9</intersection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-30,30.5,-21</points>
<intersection>-30 1</intersection>
<intersection>-21 7</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>16.5,-35,16.5,-30</points>
<intersection>-35 11</intersection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>21,-33,21,-30</points>
<intersection>-33 18</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>30.5,-21,40.5,-21</points>
<intersection>30.5 4</intersection>
<intersection>40.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>40.5,-21,40.5,-20.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>-21 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>24,-49,24,-30</points>
<intersection>-49 10</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>24,-49,41.5,-49</points>
<connection>
<GID>200</GID>
<name>IN_2</name></connection>
<intersection>24 9</intersection>
<intersection>39.5 14</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>6.5,-35,16.5,-35</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>16.5 5</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>39.5,-71.5,39.5,-49</points>
<intersection>-71.5 17</intersection>
<intersection>-64.5 16</intersection>
<intersection>-49 10</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>39.5,-64.5,42,-64.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>39.5 14</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>39.5,-71.5,42,-71.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>39.5 14</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>21,-33,23.5,-33</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>21 6</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-26,29.5,-16.5</points>
<intersection>-26 3</intersection>
<intersection>-19 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-19,29.5,-19</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-16.5,40.5,-16.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-26,40.5,-26</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection>
<intersection>39 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>39,-62.5,39,-26</points>
<intersection>-62.5 7</intersection>
<intersection>-55 8</intersection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>39,-62.5,42,-62.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>39 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>39,-55,44,-55</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>39 6</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-41,29.5,-30</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-41 3</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-30,40.5,-30</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29.5,-41,44,-41</points>
<intersection>29.5 0</intersection>
<intersection>44 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44,-41,44,-40.5</points>
<connection>
<GID>198</GID>
<name>IN_2</name></connection>
<intersection>-41 3</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-24.5,50.5,-18.5</points>
<intersection>-24.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-24.5,55,-24.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-18.5,50.5,-18.5</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-28,50.5,-26.5</points>
<intersection>-28 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-26.5,55,-26.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-28,50.5,-28</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-38.5,51,-28.5</points>
<intersection>-38.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-28.5,55,-28.5</points>
<connection>
<GID>202</GID>
<name>IN_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-38.5,51,-38.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-47,51,-30.5</points>
<intersection>-47 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-30.5,55,-30.5</points>
<connection>
<GID>202</GID>
<name>IN_3</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-47,51,-47</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-27.5,63.5,-27.5</points>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<connection>
<GID>202</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-59.5,51,-56</points>
<intersection>-59.5 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-59.5,56.5,-59.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-56,51,-56</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-63.5,51,-61.5</points>
<intersection>-63.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-61.5,56.5,-61.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-63.5,51,-63.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-70.5,51,-63.5</points>
<intersection>-70.5 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-63.5,56.5,-63.5</points>
<connection>
<GID>214</GID>
<name>IN_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-70.5,51,-70.5</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-62,63,-61.5</points>
<intersection>-62 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-62,63.5,-62</points>
<connection>
<GID>222</GID>
<name>N_in0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-61.5,63,-61.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-57,6.5,-28</points>
<intersection>-57 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-28,40.5,-28</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection>
<intersection>20.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-57,44,-57</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection>
<intersection>41.5 4</intersection>
<intersection>42 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-28,20.5,-25.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>41.5,-57,41.5,-47</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>-57 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>42,-69.5,42,-57</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-57 2</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-38.5,33.5,-18.5</points>
<intersection>-38.5 3</intersection>
<intersection>-25.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-25.5,33.5,-25.5</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-18.5,40.5,-18.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-38.5,44,-38.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>18.225,4.3,127.575,-50.975</PageViewport>
<gate>
<ID>224</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64.5,-24.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>90 </input>
<input>
<ID>IN_3</ID>91 </input>
<input>
<ID>IN_B_0</ID>87 </input>
<input>
<ID>IN_B_1</ID>86 </input>
<input>
<ID>IN_B_2</ID>85 </input>
<input>
<ID>IN_B_3</ID>84 </input>
<output>
<ID>OUT_0</ID>96 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>94 </output>
<output>
<ID>OUT_3</ID>93 </output>
<input>
<ID>carry_in</ID>97 </input>
<output>
<ID>carry_out</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_TOGGLE</type>
<position>73.5,-11.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>70.5,-11.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>67.5,-11.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>64.5,-11.5</position>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>60,-11.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_TOGGLE</type>
<position>57,-11.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_TOGGLE</type>
<position>54,-11.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_TOGGLE</type>
<position>51.5,-11.5</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>246</ID>
<type>FF_GND</type>
<position>72.5,-24.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>GA_LED</type>
<position>61,-31</position>
<input>
<ID>N_in3</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>GA_LED</type>
<position>64,-31</position>
<input>
<ID>N_in3</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>GA_LED</type>
<position>66.5,-30.5</position>
<input>
<ID>N_in3</ID>95 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>GA_LED</type>
<position>69.5,-30.5</position>
<input>
<ID>N_in3</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>GA_LED</type>
<position>52.5,-24</position>
<input>
<ID>N_in1</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>66,0</position>
<gparam>LABEL_TEXT 4 Bit Parallel Adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-20.5,64.5,-13.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>64.5,-20.5,66.5,-20.5</points>
<connection>
<GID>224</GID>
<name>IN_B_3</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-20.5,67.5,-13.5</points>
<connection>
<GID>224</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-20.5,68.5,-14.5</points>
<connection>
<GID>224</GID>
<name>IN_B_1</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-14.5,70.5,-14.5</points>
<intersection>68.5 0</intersection>
<intersection>70.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>70.5,-14.5,70.5,-13.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>73.5,-20.5,73.5,-13.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-20.5,73.5,-20.5</points>
<connection>
<GID>224</GID>
<name>IN_B_0</name></connection>
<intersection>73.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-20.5,62.5,-17</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-17 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60,-17,60,-13.5</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-17,62.5,-17</points>
<intersection>60 1</intersection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-20.5,61.5,-17.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57,-17.5,57,-13.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-17.5,61.5,-17.5</points>
<intersection>57 1</intersection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-20.5,60.5,-18.5</points>
<connection>
<GID>224</GID>
<name>IN_2</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54,-18.5,54,-13.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-18.5,60.5,-18.5</points>
<intersection>54 1</intersection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-20.5,59.5,-19.5</points>
<connection>
<GID>224</GID>
<name>IN_3</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-19.5,51.5,-13.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-19.5,59.5,-19.5</points>
<intersection>51.5 1</intersection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-30,61,-29</points>
<connection>
<GID>248</GID>
<name>N_in3</name></connection>
<intersection>-29 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>63,-29,63,-28.5</points>
<connection>
<GID>224</GID>
<name>OUT_3</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,-29,63,-29</points>
<intersection>61 0</intersection>
<intersection>63 1</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-30,64,-28.5</points>
<connection>
<GID>250</GID>
<name>N_in3</name></connection>
<connection>
<GID>224</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-29.5,66.5,-29</points>
<connection>
<GID>252</GID>
<name>N_in3</name></connection>
<intersection>-29 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>65,-29,65,-28.5</points>
<connection>
<GID>224</GID>
<name>OUT_1</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>65,-29,66.5,-29</points>
<intersection>65 1</intersection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-29.5,69.5,-29</points>
<connection>
<GID>254</GID>
<name>N_in3</name></connection>
<intersection>-29 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66,-29,66,-28.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>66,-29,69.5,-29</points>
<intersection>66 1</intersection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-23.5,72.5,-23.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<connection>
<GID>224</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-24,55,-23.5</points>
<intersection>-24 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-23.5,56.5,-23.5</points>
<connection>
<GID>224</GID>
<name>carry_out</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-24,55,-24</points>
<connection>
<GID>256</GID>
<name>N_in1</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>28.0649,-9.31351,66.4649,-28.7242</PageViewport>
<gate>
<ID>260</ID>
<type>AE_MUX_4x1</type>
<position>44.5,-21</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>100 </input>
<input>
<ID>IN_2</ID>101 </input>
<input>
<ID>IN_3</ID>102 </input>
<output>
<ID>OUT</ID>105 </output>
<input>
<ID>SEL_0</ID>104 </input>
<input>
<ID>SEL_1</ID>103 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_TOGGLE</type>
<position>37,-17</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_TOGGLE</type>
<position>37,-20</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_TOGGLE</type>
<position>37,-23</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_TOGGLE</type>
<position>37,-26</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_TOGGLE</type>
<position>43,-13</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_TOGGLE</type>
<position>47,-13</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>274</ID>
<type>GA_LED</type>
<position>51,-21</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-26,41,-24</points>
<intersection>-26 3</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-24,41.5,-24</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-26,41,-26</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-23,41,-23</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>41 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-23,41,-22</points>
<intersection>-23 1</intersection>
<intersection>-22 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41,-22,41.5,-22</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>41 3</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-20,41.5,-20</points>
<connection>
<GID>260</GID>
<name>IN_2</name></connection>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-17,41,-17</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<intersection>41 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>41,-18,41,-17</points>
<intersection>-18 6</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>41,-18,41.5,-18</points>
<connection>
<GID>260</GID>
<name>IN_3</name></connection>
<intersection>41 5</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>43,-16,43,-15</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>43,-16,44.5,-16</points>
<connection>
<GID>260</GID>
<name>SEL_1</name></connection>
<intersection>43 1</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-16,47,-15</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>45.5,-16,47,-16</points>
<connection>
<GID>260</GID>
<name>SEL_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-21,50,-21</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<connection>
<GID>274</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>-24.4098,12.3221,170.21,-86.0556</PageViewport>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>65,-7</position>
<gparam>LABEL_TEXT 8X1 MUX Using 2X1 MUX</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>AA_MUX_2x1</type>
<position>26.5,-20</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>115 </output>
<input>
<ID>SEL_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_MUX_2x1</type>
<position>26.5,-27.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>116 </output>
<input>
<ID>SEL_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_MUX_2x1</type>
<position>26.5,-35.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>117 </output>
<input>
<ID>SEL_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_MUX_2x1</type>
<position>26.5,-44</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>118 </output>
<input>
<ID>SEL_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_MUX_2x1</type>
<position>40,-23.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>119 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_MUX_2x1</type>
<position>40,-39</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>120 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_MUX_2x1</type>
<position>53,-29</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>123 </output>
<input>
<ID>SEL_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_TOGGLE</type>
<position>20,-19</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_TOGGLE</type>
<position>20,-21.5</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_TOGGLE</type>
<position>20,-26</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_TOGGLE</type>
<position>20,-29</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_TOGGLE</type>
<position>20,-33.5</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_TOGGLE</type>
<position>20,-37</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_TOGGLE</type>
<position>20,-42</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_TOGGLE</type>
<position>20,-45</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_TOGGLE</type>
<position>17,-12</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_TOGGLE</type>
<position>39.5,-17</position>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_TOGGLE</type>
<position>53,-21</position>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>314</ID>
<type>GA_LED</type>
<position>57.5,-29</position>
<input>
<ID>N_in0</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-43,23,-42</points>
<intersection>-43 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-43,24.5,-43</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-42,23,-42</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-45,24.5,-45</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-34.5,23,-33.5</points>
<intersection>-34.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-34.5,24.5,-34.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-33.5,23,-33.5</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-37,23.5,-36.5</points>
<intersection>-37 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-36.5,24.5,-36.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-37,23.5,-37</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-26.5,23,-26</points>
<intersection>-26.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-26.5,24.5,-26.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-26,23,-26</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-29,23,-28.5</points>
<intersection>-29 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-28.5,24.5,-28.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-29,23,-29</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-19,24.5,-19</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-19,24.5,-19</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-21.5,23,-21</points>
<intersection>-21.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-21,24.5,-21</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-21.5,23,-21.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-40,17,-14</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<intersection>-40 12</intersection>
<intersection>-31.5 13</intersection>
<intersection>-24.5 7</intersection>
<intersection>-17.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>17,-24.5,26.5,-24.5</points>
<intersection>17 0</intersection>
<intersection>26.5 15</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17,-17.5,26.5,-17.5</points>
<connection>
<GID>278</GID>
<name>SEL_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>17,-40,26.5,-40</points>
<intersection>17 0</intersection>
<intersection>26.5 16</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>17,-31.5,26.5,-31.5</points>
<intersection>17 0</intersection>
<intersection>26.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>26.5,-33,26.5,-31.5</points>
<connection>
<GID>282</GID>
<name>SEL_0</name></connection>
<intersection>-31.5 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>26.5,-25,26.5,-24.5</points>
<connection>
<GID>280</GID>
<name>SEL_0</name></connection>
<intersection>-24.5 7</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>26.5,-41.5,26.5,-40</points>
<connection>
<GID>284</GID>
<name>SEL_0</name></connection>
<intersection>-40 12</intersection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-22.5,32.5,-20</points>
<intersection>-22.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-22.5,38,-22.5</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-20,32.5,-20</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-27.5,32.5,-24.5</points>
<intersection>-27.5 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-24.5,38,-24.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-27.5,32.5,-27.5</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-38,32.5,-35.5</points>
<intersection>-38 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-38,38,-38</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-35.5,32.5,-35.5</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-44,32.5,-40</points>
<intersection>-44 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-40,38,-40</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-44,32.5,-44</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-28,46.5,-23.5</points>
<intersection>-28 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-28,51,-28</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-23.5,46.5,-23.5</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-39,46.5,-30</points>
<intersection>-39 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-30,51,-30</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-39,46.5,-39</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-36.5,43.5,-20</points>
<intersection>-36.5 4</intersection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39.5,-20,39.5,-19</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-20,43.5,-20</points>
<intersection>39.5 1</intersection>
<intersection>40 6</intersection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40,-36.5,43.5,-36.5</points>
<connection>
<GID>288</GID>
<name>SEL_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-21,40,-20</points>
<connection>
<GID>286</GID>
<name>SEL_0</name></connection>
<intersection>-20 2</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-26.5,53,-23</points>
<connection>
<GID>290</GID>
<name>SEL_0</name></connection>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-29,56.5,-29</points>
<connection>
<GID>314</GID>
<name>N_in0</name></connection>
<connection>
<GID>290</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>