<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>501.616,517.939,603.501,467.579</PageViewport>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>556,506.5</position>
<gparam>LABEL_TEXT 4 bit synchronous up counter using T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BE_JKFF_LOW</type>
<position>526.5,492</position>
<input>
<ID>J</ID>16 </input>
<input>
<ID>K</ID>16 </input>
<output>
<ID>Q</ID>7 </output>
<input>
<ID>clock</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>BE_JKFF_LOW</type>
<position>534.5,490.5</position>
<input>
<ID>J</ID>7 </input>
<input>
<ID>K</ID>7 </input>
<output>
<ID>Q</ID>12 </output>
<input>
<ID>clock</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>18</ID>
<type>BE_JKFF_LOW</type>
<position>547.5,492</position>
<input>
<ID>J</ID>8 </input>
<input>
<ID>K</ID>8 </input>
<output>
<ID>Q</ID>13 </output>
<input>
<ID>clock</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>BE_JKFF_LOW</type>
<position>565.5,492</position>
<input>
<ID>J</ID>9 </input>
<input>
<ID>K</ID>9 </input>
<output>
<ID>Q</ID>15 </output>
<input>
<ID>clock</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>22</ID>
<type>BB_CLOCK</type>
<position>515,492</position>
<output>
<ID>CLK</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>541.5,499</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>556.5,499</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>587.5,493</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>15 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>520,490</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,479.5,530,492.5</points>
<intersection>479.5 7</intersection>
<intersection>488.5 12</intersection>
<intersection>492.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529.5,492.5,531.5,492.5</points>
<connection>
<GID>16</GID>
<name>J</name></connection>
<intersection>529.5 11</intersection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>530,479.5,581.5,479.5</points>
<intersection>530 0</intersection>
<intersection>538.5 9</intersection>
<intersection>581.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>581.5,479.5,581.5,492</points>
<intersection>479.5 7</intersection>
<intersection>492 10</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>538.5,479.5,538.5,500</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>479.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>581.5,492,584.5,492</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>581.5 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>529.5,492.5,529.5,494</points>
<connection>
<GID>14</GID>
<name>Q</name></connection>
<intersection>492.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>530,488.5,531.5,488.5</points>
<connection>
<GID>16</GID>
<name>K</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543.5,490,543.5,500</points>
<intersection>490 2</intersection>
<intersection>494 1</intersection>
<intersection>499 6</intersection>
<intersection>500 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>543.5,494,544.5,494</points>
<connection>
<GID>18</GID>
<name>J</name></connection>
<intersection>543.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>543.5,490,544.5,490</points>
<connection>
<GID>18</GID>
<name>K</name></connection>
<intersection>543.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>543.5,500,553.5,500</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>543.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>543.5,499,544.5,499</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>543.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>560,490,560,499</points>
<intersection>490 2</intersection>
<intersection>494 1</intersection>
<intersection>499 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>560,494,562.5,494</points>
<connection>
<GID>20</GID>
<name>J</name></connection>
<intersection>560 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>560,490,562.5,490</points>
<connection>
<GID>20</GID>
<name>K</name></connection>
<intersection>560 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>559.5,499,560,499</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>560 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537.5,484,537.5,498</points>
<connection>
<GID>16</GID>
<name>Q</name></connection>
<intersection>484 3</intersection>
<intersection>498 8</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>537.5,484,580,484</points>
<intersection>537.5 0</intersection>
<intersection>580 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>580,484,580,493</points>
<intersection>484 3</intersection>
<intersection>493 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>580,493,584.5,493</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>580 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>537.5,498,538.5,498</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>537.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>552,487.5,552,493</points>
<intersection>487.5 1</intersection>
<intersection>493 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>552,487.5,579.5,487.5</points>
<intersection>552 0</intersection>
<intersection>553.5 6</intersection>
<intersection>579.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>550.5,493,552,493</points>
<intersection>550.5 3</intersection>
<intersection>552 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>550.5,493,550.5,494</points>
<connection>
<GID>18</GID>
<name>Q</name></connection>
<intersection>493 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>579.5,487.5,579.5,494</points>
<intersection>487.5 1</intersection>
<intersection>494 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>579.5,494,584.5,494</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<intersection>579.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>553.5,487.5,553.5,498</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>487.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,502,561.5,502</points>
<intersection>519 6</intersection>
<intersection>522.5 5</intersection>
<intersection>531.5 4</intersection>
<intersection>544.5 8</intersection>
<intersection>561.5 10</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>531.5,490.5,531.5,502</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>502 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>522.5,492,522.5,502</points>
<intersection>492 12</intersection>
<intersection>502 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>519,492,519,502</points>
<connection>
<GID>22</GID>
<name>CLK</name></connection>
<intersection>502 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>544.5,492,544.5,502</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>502 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>561.5,492,561.5,502</points>
<intersection>492 11</intersection>
<intersection>502 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>561.5,492,562.5,492</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<intersection>561.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>522.5,492,523.5,492</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>522.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>568.5,495,584.5,495</points>
<connection>
<GID>34</GID>
<name>IN_3</name></connection>
<intersection>568.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>568.5,494,568.5,495</points>
<connection>
<GID>20</GID>
<name>Q</name></connection>
<intersection>495 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>523.5,490,523.5,494</points>
<connection>
<GID>14</GID>
<name>K</name></connection>
<connection>
<GID>14</GID>
<name>J</name></connection>
<intersection>490 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>522,490,523.5,490</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>523.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-12,-3,110.4,-63.5</PageViewport>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>46,-5</position>
<gparam>LABEL_TEXT 0-2-3-6-4-0 using D flipflop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AE_DFF_LOW</type>
<position>24,-26.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUTINV_0</ID>19 </output>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_DFF_LOW</type>
<position>42,-26.5</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>18 </output>
<input>
<ID>clock</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_DFF_LOW</type>
<position>56.5,-30.5</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUTINV_0</ID>26 </output>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND3</type>
<position>8,-16.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>50</ID>
<type>BB_CLOCK</type>
<position>8,-27.5</position>
<output>
<ID>CLK</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 12</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>51,-13.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR2</type>
<position>67,-18</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>88,-39.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>23 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-10.5,47,-10.5</points>
<intersection>4 4</intersection>
<intersection>47 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,-39.5,47,-10.5</points>
<intersection>-39.5 7</intersection>
<intersection>-24.5 8</intersection>
<intersection>-14.5 6</intersection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>4,-16.5,4,-10.5</points>
<intersection>-16.5 5</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4,-16.5,5,-16.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>4 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47,-14.5,48,-14.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>47 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>47,-39.5,85,-39.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>47 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>45,-24.5,47,-24.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>47 3</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-38.5,2.5,-18.5</points>
<intersection>-38.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-18.5,5,-18.5</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-38.5,27,-38.5</points>
<intersection>2.5 0</intersection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-38.5,27,-27.5</points>
<connection>
<GID>40</GID>
<name>OUTINV_0</name></connection>
<intersection>-38.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-24.5,16,-16.5</points>
<intersection>-24.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-24.5,21,-24.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-16.5,16,-16.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-43,52,-43</points>
<intersection>12 6</intersection>
<intersection>21 5</intersection>
<intersection>35.5 4</intersection>
<intersection>52 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>35.5,-43,35.5,-27.5</points>
<intersection>-43 1</intersection>
<intersection>-27.5 10</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>21,-43,21,-27.5</points>
<connection>
<GID>40</GID>
<name>clock</name></connection>
<intersection>-43 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>12,-43,12,-27.5</points>
<connection>
<GID>50</GID>
<name>CLK</name></connection>
<intersection>-43 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>52,-43,52,-31.5</points>
<intersection>-43 1</intersection>
<intersection>-31.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>52,-31.5,53.5,-31.5</points>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<intersection>52 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>35.5,-27.5,39,-27.5</points>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<intersection>35.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-55,29.5,-24.5</points>
<intersection>-55 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-55,72,-55</points>
<intersection>29.5 0</intersection>
<intersection>64 6</intersection>
<intersection>72 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-24.5,29.5,-24.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72,-55,72,-40.5</points>
<intersection>-55 1</intersection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>72,-40.5,85,-40.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>72 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64,-55,64,-17</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-25.5,48,-12.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48,-25.5,62,-25.5</points>
<intersection>48 0</intersection>
<intersection>62 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62,-38.5,62,-25.5</points>
<intersection>-38.5 4</intersection>
<intersection>-28.5 5</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,-38.5,85,-38.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>62 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59.5,-28.5,62,-28.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>62 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-19,59,-13.5</points>
<intersection>-19 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-19,64,-19</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-13.5,59,-13.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-24,61.5,-22</points>
<intersection>-24 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-22,61.5,-22</points>
<intersection>53.5 4</intersection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-24,70,-24</points>
<intersection>61.5 0</intersection>
<intersection>70 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70,-24,70,-18</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-28.5,53.5,-22</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-18.5,49,-13</points>
<intersection>-18.5 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-13,49,-13</points>
<intersection>5 7</intersection>
<intersection>33 4</intersection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-18.5,60.5,-18.5</points>
<intersection>49 0</intersection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-31.5,60.5,-18.5</points>
<intersection>-31.5 5</intersection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>33,-24.5,33,-13</points>
<intersection>-24.5 6</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>59.5,-31.5,60.5,-31.5</points>
<connection>
<GID>44</GID>
<name>OUTINV_0</name></connection>
<intersection>60.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>33,-24.5,39,-24.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>33 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>5,-14.5,5,-13</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>